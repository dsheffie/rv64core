`include "machine.vh"
module ppa32(A, B, Y);
   input [31:0] A;
   input [31:0] B;
   output [31:0] Y;
`ifdef FPGA
   assign Y = A+B;
`else
   wire 	 pp_0 = A[0] ^ B[0];
   wire 	 gg_0 = A[0] & B[0];
   wire 	 pp_1 = A[1] ^ B[1];
   wire 	 gg_1 = A[1] & B[1];
   wire 	 pp_2 = A[2] ^ B[2];
   wire 	 gg_2 = A[2] & B[2];
   wire 	 pp_3 = A[3] ^ B[3];
   wire 	 gg_3 = A[3] & B[3];
   wire 	 pp_4 = A[4] ^ B[4];
   wire 	 gg_4 = A[4] & B[4];
   wire 	 pp_5 = A[5] ^ B[5];
   wire 	 gg_5 = A[5] & B[5];
   wire 	 pp_6 = A[6] ^ B[6];
   wire 	 gg_6 = A[6] & B[6];
   wire 	 pp_7 = A[7] ^ B[7];
   wire 	 gg_7 = A[7] & B[7];
   wire 	 pp_8 = A[8] ^ B[8];
   wire 	 gg_8 = A[8] & B[8];
   wire 	 pp_9 = A[9] ^ B[9];
   wire 	 gg_9 = A[9] & B[9];
   wire 	 pp_10 = A[10] ^ B[10];
   wire 	 gg_10 = A[10] & B[10];
   wire 	 pp_11 = A[11] ^ B[11];
   wire 	 gg_11 = A[11] & B[11];
   wire 	 pp_12 = A[12] ^ B[12];
   wire 	 gg_12 = A[12] & B[12];
   wire 	 pp_13 = A[13] ^ B[13];
   wire 	 gg_13 = A[13] & B[13];
   wire 	 pp_14 = A[14] ^ B[14];
   wire 	 gg_14 = A[14] & B[14];
   wire 	 pp_15 = A[15] ^ B[15];
   wire 	 gg_15 = A[15] & B[15];
   wire 	 pp_16 = A[16] ^ B[16];
   wire 	 gg_16 = A[16] & B[16];
   wire 	 pp_17 = A[17] ^ B[17];
   wire 	 gg_17 = A[17] & B[17];
   wire 	 pp_18 = A[18] ^ B[18];
   wire 	 gg_18 = A[18] & B[18];
   wire 	 pp_19 = A[19] ^ B[19];
   wire 	 gg_19 = A[19] & B[19];
   wire 	 pp_20 = A[20] ^ B[20];
   wire 	 gg_20 = A[20] & B[20];
   wire 	 pp_21 = A[21] ^ B[21];
   wire 	 gg_21 = A[21] & B[21];
   wire 	 pp_22 = A[22] ^ B[22];
   wire 	 gg_22 = A[22] & B[22];
   wire 	 pp_23 = A[23] ^ B[23];
   wire 	 gg_23 = A[23] & B[23];
   wire 	 pp_24 = A[24] ^ B[24];
   wire 	 gg_24 = A[24] & B[24];
   wire 	 pp_25 = A[25] ^ B[25];
   wire 	 gg_25 = A[25] & B[25];
   wire 	 pp_26 = A[26] ^ B[26];
   wire 	 gg_26 = A[26] & B[26];
   wire 	 pp_27 = A[27] ^ B[27];
   wire 	 gg_27 = A[27] & B[27];
   wire 	 pp_28 = A[28] ^ B[28];
   wire 	 gg_28 = A[28] & B[28];
   wire 	 pp_29 = A[29] ^ B[29];
   wire 	 gg_29 = A[29] & B[29];
   wire 	 pp_30 = A[30] ^ B[30];
   wire 	 gg_30 = A[30] & B[30];
   wire 	 pp_31 = A[31] ^ B[31];
   wire 	 gg_31 = A[31] & B[31];
   wire 	 pp_1_pp_0 = pp_1 & pp_0;
   wire 	 gg_1_gg_0 = (gg_0 & pp_1) | gg_1;
   wire 	 pp_2_pp_1 = pp_2 & pp_1;
   wire 	 gg_2_gg_1 = (gg_1 & pp_2) | gg_2;
   wire 	 pp_3_pp_2 = pp_3 & pp_2;
   wire 	 gg_3_gg_2 = (gg_2 & pp_3) | gg_3;
   wire 	 pp_4_pp_3 = pp_4 & pp_3;
   wire 	 gg_4_gg_3 = (gg_3 & pp_4) | gg_4;
   wire 	 pp_5_pp_4 = pp_5 & pp_4;
   wire 	 gg_5_gg_4 = (gg_4 & pp_5) | gg_5;
   wire 	 pp_6_pp_5 = pp_6 & pp_5;
   wire 	 gg_6_gg_5 = (gg_5 & pp_6) | gg_6;
   wire 	 pp_7_pp_6 = pp_7 & pp_6;
   wire 	 gg_7_gg_6 = (gg_6 & pp_7) | gg_7;
   wire 	 pp_8_pp_7 = pp_8 & pp_7;
   wire 	 gg_8_gg_7 = (gg_7 & pp_8) | gg_8;
   wire 	 pp_9_pp_8 = pp_9 & pp_8;
   wire 	 gg_9_gg_8 = (gg_8 & pp_9) | gg_9;
   wire 	 pp_10_pp_9 = pp_10 & pp_9;
   wire 	 gg_10_gg_9 = (gg_9 & pp_10) | gg_10;
   wire 	 pp_11_pp_10 = pp_11 & pp_10;
   wire 	 gg_11_gg_10 = (gg_10 & pp_11) | gg_11;
   wire 	 pp_12_pp_11 = pp_12 & pp_11;
   wire 	 gg_12_gg_11 = (gg_11 & pp_12) | gg_12;
   wire 	 pp_13_pp_12 = pp_13 & pp_12;
   wire 	 gg_13_gg_12 = (gg_12 & pp_13) | gg_13;
   wire 	 pp_14_pp_13 = pp_14 & pp_13;
   wire 	 gg_14_gg_13 = (gg_13 & pp_14) | gg_14;
   wire 	 pp_15_pp_14 = pp_15 & pp_14;
   wire 	 gg_15_gg_14 = (gg_14 & pp_15) | gg_15;
   wire 	 pp_16_pp_15 = pp_16 & pp_15;
   wire 	 gg_16_gg_15 = (gg_15 & pp_16) | gg_16;
   wire 	 pp_17_pp_16 = pp_17 & pp_16;
   wire 	 gg_17_gg_16 = (gg_16 & pp_17) | gg_17;
   wire 	 pp_18_pp_17 = pp_18 & pp_17;
   wire 	 gg_18_gg_17 = (gg_17 & pp_18) | gg_18;
   wire 	 pp_19_pp_18 = pp_19 & pp_18;
   wire 	 gg_19_gg_18 = (gg_18 & pp_19) | gg_19;
   wire 	 pp_20_pp_19 = pp_20 & pp_19;
   wire 	 gg_20_gg_19 = (gg_19 & pp_20) | gg_20;
   wire 	 pp_21_pp_20 = pp_21 & pp_20;
   wire 	 gg_21_gg_20 = (gg_20 & pp_21) | gg_21;
   wire 	 pp_22_pp_21 = pp_22 & pp_21;
   wire 	 gg_22_gg_21 = (gg_21 & pp_22) | gg_22;
   wire 	 pp_23_pp_22 = pp_23 & pp_22;
   wire 	 gg_23_gg_22 = (gg_22 & pp_23) | gg_23;
   wire 	 pp_24_pp_23 = pp_24 & pp_23;
   wire 	 gg_24_gg_23 = (gg_23 & pp_24) | gg_24;
   wire 	 pp_25_pp_24 = pp_25 & pp_24;
   wire 	 gg_25_gg_24 = (gg_24 & pp_25) | gg_25;
   wire 	 pp_26_pp_25 = pp_26 & pp_25;
   wire 	 gg_26_gg_25 = (gg_25 & pp_26) | gg_26;
   wire 	 pp_27_pp_26 = pp_27 & pp_26;
   wire 	 gg_27_gg_26 = (gg_26 & pp_27) | gg_27;
   wire 	 pp_28_pp_27 = pp_28 & pp_27;
   wire 	 gg_28_gg_27 = (gg_27 & pp_28) | gg_28;
   wire 	 pp_29_pp_28 = pp_29 & pp_28;
   wire 	 gg_29_gg_28 = (gg_28 & pp_29) | gg_29;
   wire 	 pp_30_pp_29 = pp_30 & pp_29;
   wire 	 gg_30_gg_29 = (gg_29 & pp_30) | gg_30;
   wire 	 pp_31_pp_30 = pp_31 & pp_30;
   wire 	 gg_31_gg_30 = (gg_30 & pp_31) | gg_31;
   wire 	 pp_2_pp_1_pp_0 = pp_2_pp_1 & pp_0;
   wire 	 gg_2_gg_1_gg_0 = (gg_0 & pp_2_pp_1) | gg_2_gg_1;
   wire 	 pp_3_pp_2_pp_1_pp_0 = pp_3_pp_2 & pp_1_pp_0;
   wire 	 gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_3_pp_2) | gg_3_gg_2;
   wire 	 pp_4_pp_3_pp_2_pp_1 = pp_4_pp_3 & pp_2_pp_1;
   wire 	 gg_4_gg_3_gg_2_gg_1 = (gg_2_gg_1 & pp_4_pp_3) | gg_4_gg_3;
   wire 	 pp_5_pp_4_pp_3_pp_2 = pp_5_pp_4 & pp_3_pp_2;
   wire 	 gg_5_gg_4_gg_3_gg_2 = (gg_3_gg_2 & pp_5_pp_4) | gg_5_gg_4;
   wire 	 pp_6_pp_5_pp_4_pp_3 = pp_6_pp_5 & pp_4_pp_3;
   wire 	 gg_6_gg_5_gg_4_gg_3 = (gg_4_gg_3 & pp_6_pp_5) | gg_6_gg_5;
   wire 	 pp_7_pp_6_pp_5_pp_4 = pp_7_pp_6 & pp_5_pp_4;
   wire 	 gg_7_gg_6_gg_5_gg_4 = (gg_5_gg_4 & pp_7_pp_6) | gg_7_gg_6;
   wire 	 pp_8_pp_7_pp_6_pp_5 = pp_8_pp_7 & pp_6_pp_5;
   wire 	 gg_8_gg_7_gg_6_gg_5 = (gg_6_gg_5 & pp_8_pp_7) | gg_8_gg_7;
   wire 	 pp_9_pp_8_pp_7_pp_6 = pp_9_pp_8 & pp_7_pp_6;
   wire 	 gg_9_gg_8_gg_7_gg_6 = (gg_7_gg_6 & pp_9_pp_8) | gg_9_gg_8;
   wire 	 pp_10_pp_9_pp_8_pp_7 = pp_10_pp_9 & pp_8_pp_7;
   wire 	 gg_10_gg_9_gg_8_gg_7 = (gg_8_gg_7 & pp_10_pp_9) | gg_10_gg_9;
   wire 	 pp_11_pp_10_pp_9_pp_8 = pp_11_pp_10 & pp_9_pp_8;
   wire 	 gg_11_gg_10_gg_9_gg_8 = (gg_9_gg_8 & pp_11_pp_10) | gg_11_gg_10;
   wire 	 pp_12_pp_11_pp_10_pp_9 = pp_12_pp_11 & pp_10_pp_9;
   wire 	 gg_12_gg_11_gg_10_gg_9 = (gg_10_gg_9 & pp_12_pp_11) | gg_12_gg_11;
   wire 	 pp_13_pp_12_pp_11_pp_10 = pp_13_pp_12 & pp_11_pp_10;
   wire 	 gg_13_gg_12_gg_11_gg_10 = (gg_11_gg_10 & pp_13_pp_12) | gg_13_gg_12;
   wire 	 pp_14_pp_13_pp_12_pp_11 = pp_14_pp_13 & pp_12_pp_11;
   wire 	 gg_14_gg_13_gg_12_gg_11 = (gg_12_gg_11 & pp_14_pp_13) | gg_14_gg_13;
   wire 	 pp_15_pp_14_pp_13_pp_12 = pp_15_pp_14 & pp_13_pp_12;
   wire 	 gg_15_gg_14_gg_13_gg_12 = (gg_13_gg_12 & pp_15_pp_14) | gg_15_gg_14;
   wire 	 pp_16_pp_15_pp_14_pp_13 = pp_16_pp_15 & pp_14_pp_13;
   wire 	 gg_16_gg_15_gg_14_gg_13 = (gg_14_gg_13 & pp_16_pp_15) | gg_16_gg_15;
   wire 	 pp_17_pp_16_pp_15_pp_14 = pp_17_pp_16 & pp_15_pp_14;
   wire 	 gg_17_gg_16_gg_15_gg_14 = (gg_15_gg_14 & pp_17_pp_16) | gg_17_gg_16;
   wire 	 pp_18_pp_17_pp_16_pp_15 = pp_18_pp_17 & pp_16_pp_15;
   wire 	 gg_18_gg_17_gg_16_gg_15 = (gg_16_gg_15 & pp_18_pp_17) | gg_18_gg_17;
   wire 	 pp_19_pp_18_pp_17_pp_16 = pp_19_pp_18 & pp_17_pp_16;
   wire 	 gg_19_gg_18_gg_17_gg_16 = (gg_17_gg_16 & pp_19_pp_18) | gg_19_gg_18;
   wire 	 pp_20_pp_19_pp_18_pp_17 = pp_20_pp_19 & pp_18_pp_17;
   wire 	 gg_20_gg_19_gg_18_gg_17 = (gg_18_gg_17 & pp_20_pp_19) | gg_20_gg_19;
   wire 	 pp_21_pp_20_pp_19_pp_18 = pp_21_pp_20 & pp_19_pp_18;
   wire 	 gg_21_gg_20_gg_19_gg_18 = (gg_19_gg_18 & pp_21_pp_20) | gg_21_gg_20;
   wire 	 pp_22_pp_21_pp_20_pp_19 = pp_22_pp_21 & pp_20_pp_19;
   wire 	 gg_22_gg_21_gg_20_gg_19 = (gg_20_gg_19 & pp_22_pp_21) | gg_22_gg_21;
   wire 	 pp_23_pp_22_pp_21_pp_20 = pp_23_pp_22 & pp_21_pp_20;
   wire 	 gg_23_gg_22_gg_21_gg_20 = (gg_21_gg_20 & pp_23_pp_22) | gg_23_gg_22;
   wire 	 pp_24_pp_23_pp_22_pp_21 = pp_24_pp_23 & pp_22_pp_21;
   wire 	 gg_24_gg_23_gg_22_gg_21 = (gg_22_gg_21 & pp_24_pp_23) | gg_24_gg_23;
   wire 	 pp_25_pp_24_pp_23_pp_22 = pp_25_pp_24 & pp_23_pp_22;
   wire 	 gg_25_gg_24_gg_23_gg_22 = (gg_23_gg_22 & pp_25_pp_24) | gg_25_gg_24;
   wire 	 pp_26_pp_25_pp_24_pp_23 = pp_26_pp_25 & pp_24_pp_23;
   wire 	 gg_26_gg_25_gg_24_gg_23 = (gg_24_gg_23 & pp_26_pp_25) | gg_26_gg_25;
   wire 	 pp_27_pp_26_pp_25_pp_24 = pp_27_pp_26 & pp_25_pp_24;
   wire 	 gg_27_gg_26_gg_25_gg_24 = (gg_25_gg_24 & pp_27_pp_26) | gg_27_gg_26;
   wire 	 pp_28_pp_27_pp_26_pp_25 = pp_28_pp_27 & pp_26_pp_25;
   wire 	 gg_28_gg_27_gg_26_gg_25 = (gg_26_gg_25 & pp_28_pp_27) | gg_28_gg_27;
   wire 	 pp_29_pp_28_pp_27_pp_26 = pp_29_pp_28 & pp_27_pp_26;
   wire 	 gg_29_gg_28_gg_27_gg_26 = (gg_27_gg_26 & pp_29_pp_28) | gg_29_gg_28;
   wire 	 pp_30_pp_29_pp_28_pp_27 = pp_30_pp_29 & pp_28_pp_27;
   wire 	 gg_30_gg_29_gg_28_gg_27 = (gg_28_gg_27 & pp_30_pp_29) | gg_30_gg_29;
   wire 	 pp_31_pp_30_pp_29_pp_28 = pp_31_pp_30 & pp_29_pp_28;
   wire 	 gg_31_gg_30_gg_29_gg_28 = (gg_29_gg_28 & pp_31_pp_30) | gg_31_gg_30;
   wire 	 pp_4_pp_3_pp_2_pp_1_pp_0 = pp_4_pp_3_pp_2_pp_1 & pp_0;
   wire 	 gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_4_pp_3_pp_2_pp_1) | gg_4_gg_3_gg_2_gg_1;
   wire 	 pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
   wire 	 gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_5_pp_4_pp_3_pp_2) | gg_5_gg_4_gg_3_gg_2;
   wire 	 pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
   wire 	 gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_6_pp_5_pp_4_pp_3) | gg_6_gg_5_gg_4_gg_3;
   wire 	 pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_7_pp_6_pp_5_pp_4) | gg_7_gg_6_gg_5_gg_4;
   wire 	 pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 = pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1;
   wire 	 gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 = (gg_4_gg_3_gg_2_gg_1 & pp_8_pp_7_pp_6_pp_5) | gg_8_gg_7_gg_6_gg_5;
   wire 	 pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 = pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2;
   wire 	 gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 = (gg_5_gg_4_gg_3_gg_2 & pp_9_pp_8_pp_7_pp_6) | gg_9_gg_8_gg_7_gg_6;
   wire 	 pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 = pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3;
   wire 	 gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 = (gg_6_gg_5_gg_4_gg_3 & pp_10_pp_9_pp_8_pp_7) | gg_10_gg_9_gg_8_gg_7;
   wire 	 pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 = pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4;
   wire 	 gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 = (gg_7_gg_6_gg_5_gg_4 & pp_11_pp_10_pp_9_pp_8) | gg_11_gg_10_gg_9_gg_8;
   wire 	 pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 = pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5;
   wire 	 gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 = (gg_8_gg_7_gg_6_gg_5 & pp_12_pp_11_pp_10_pp_9) | gg_12_gg_11_gg_10_gg_9;
   wire 	 pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 = pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6;
   wire 	 gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 = (gg_9_gg_8_gg_7_gg_6 & pp_13_pp_12_pp_11_pp_10) | gg_13_gg_12_gg_11_gg_10;
   wire 	 pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 = pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7;
   wire 	 gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 = (gg_10_gg_9_gg_8_gg_7 & pp_14_pp_13_pp_12_pp_11) | gg_14_gg_13_gg_12_gg_11;
   wire 	 pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 = pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8;
   wire 	 gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 = (gg_11_gg_10_gg_9_gg_8 & pp_15_pp_14_pp_13_pp_12) | gg_15_gg_14_gg_13_gg_12;
   wire 	 pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 = pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9;
   wire 	 gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 = (gg_12_gg_11_gg_10_gg_9 & pp_16_pp_15_pp_14_pp_13) | gg_16_gg_15_gg_14_gg_13;
   wire 	 pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 = pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10;
   wire 	 gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 = (gg_13_gg_12_gg_11_gg_10 & pp_17_pp_16_pp_15_pp_14) | gg_17_gg_16_gg_15_gg_14;
   wire 	 pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 = pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11;
   wire 	 gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 = (gg_14_gg_13_gg_12_gg_11 & pp_18_pp_17_pp_16_pp_15) | gg_18_gg_17_gg_16_gg_15;
   wire 	 pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 = pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12;
   wire 	 gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 = (gg_15_gg_14_gg_13_gg_12 & pp_19_pp_18_pp_17_pp_16) | gg_19_gg_18_gg_17_gg_16;
   wire 	 pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 = pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13;
   wire 	 gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 = (gg_16_gg_15_gg_14_gg_13 & pp_20_pp_19_pp_18_pp_17) | gg_20_gg_19_gg_18_gg_17;
   wire 	 pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 = pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14;
   wire 	 gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 = (gg_17_gg_16_gg_15_gg_14 & pp_21_pp_20_pp_19_pp_18) | gg_21_gg_20_gg_19_gg_18;
   wire 	 pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 = pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15;
   wire 	 gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 = (gg_18_gg_17_gg_16_gg_15 & pp_22_pp_21_pp_20_pp_19) | gg_22_gg_21_gg_20_gg_19;
   wire 	 pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 = pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16;
   wire 	 gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 = (gg_19_gg_18_gg_17_gg_16 & pp_23_pp_22_pp_21_pp_20) | gg_23_gg_22_gg_21_gg_20;
   wire 	 pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 = pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17;
   wire 	 gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 = (gg_20_gg_19_gg_18_gg_17 & pp_24_pp_23_pp_22_pp_21) | gg_24_gg_23_gg_22_gg_21;
   wire 	 pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 = pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18;
   wire 	 gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 = (gg_21_gg_20_gg_19_gg_18 & pp_25_pp_24_pp_23_pp_22) | gg_25_gg_24_gg_23_gg_22;
   wire 	 pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 = pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19;
   wire 	 gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 = (gg_22_gg_21_gg_20_gg_19 & pp_26_pp_25_pp_24_pp_23) | gg_26_gg_25_gg_24_gg_23;
   wire 	 pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 = pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20;
   wire 	 gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 = (gg_23_gg_22_gg_21_gg_20 & pp_27_pp_26_pp_25_pp_24) | gg_27_gg_26_gg_25_gg_24;
   wire 	 pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 = pp_28_pp_27_pp_26_pp_25 & pp_24_pp_23_pp_22_pp_21;
   wire 	 gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 = (gg_24_gg_23_gg_22_gg_21 & pp_28_pp_27_pp_26_pp_25) | gg_28_gg_27_gg_26_gg_25;
   wire 	 pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 = pp_29_pp_28_pp_27_pp_26 & pp_25_pp_24_pp_23_pp_22;
   wire 	 gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 = (gg_25_gg_24_gg_23_gg_22 & pp_29_pp_28_pp_27_pp_26) | gg_29_gg_28_gg_27_gg_26;
   wire 	 pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 = pp_30_pp_29_pp_28_pp_27 & pp_26_pp_25_pp_24_pp_23;
   wire 	 gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 = (gg_26_gg_25_gg_24_gg_23 & pp_30_pp_29_pp_28_pp_27) | gg_30_gg_29_gg_28_gg_27;
   wire 	 pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 = pp_31_pp_30_pp_29_pp_28 & pp_27_pp_26_pp_25_pp_24;
   wire 	 gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 = (gg_27_gg_26_gg_25_gg_24 & pp_31_pp_30_pp_29_pp_28) | gg_31_gg_30_gg_29_gg_28;
   wire 	 pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 & pp_0;
   wire 	 gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1) | gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1;
   wire 	 pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
   wire 	 gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2) | gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2;
   wire 	 pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
   wire 	 gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3) | gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3;
   wire 	 pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4) | gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4;
   wire 	 pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_4_gg_3_gg_2_gg_1_gg_0 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5) | gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5;
   wire 	 pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6) | gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6;
   wire 	 pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7) | gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7;
   wire 	 pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8) | gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8;
   wire 	 pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 = pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1;
   wire 	 gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 = (gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9) | gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9;
   wire 	 pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 = pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2;
   wire 	 gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 = (gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10) | gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10;
   wire 	 pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 = pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3;
   wire 	 gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 = (gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11) | gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11;
   wire 	 pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 = pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4;
   wire 	 gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 = (gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12) | gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12;
   wire 	 pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 = pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5;
   wire 	 gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 = (gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13) | gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13;
   wire 	 pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 = pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6;
   wire 	 gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 = (gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14) | gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14;
   wire 	 pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 = pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7;
   wire 	 gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 = (gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15) | gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15;
   wire 	 pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 = pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8;
   wire 	 gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 = (gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16) | gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16;
   wire 	 pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 = pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9;
   wire 	 gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 = (gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17) | gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17;
   wire 	 pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 = pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10;
   wire 	 gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 = (gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18) | gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18;
   wire 	 pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 = pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11;
   wire 	 gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 = (gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19) | gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19;
   wire 	 pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 = pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12;
   wire 	 gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 = (gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20) | gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20;
   wire 	 pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 = pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13;
   wire 	 gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 = (gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21) | gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21;
   wire 	 pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 = pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14;
   wire 	 gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 = (gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22) | gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22;
   wire 	 pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 = pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15;
   wire 	 gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 = (gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23) | gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23;
   wire 	 pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 = pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16;
   wire 	 gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 = (gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24) | gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24;
   wire 	 pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 & pp_0;
   wire 	 gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1) | gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1;
   wire 	 pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
   wire 	 gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2) | gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2;
   wire 	 pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
   wire 	 gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3) | gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3;
   wire 	 pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4) | gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4;
   wire 	 pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_4_gg_3_gg_2_gg_1_gg_0 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5) | gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5;
   wire 	 pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6) | gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6;
   wire 	 pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7) | gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7;
   wire 	 pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8) | gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8;
   wire 	 pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9) | gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9;
   wire 	 pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10) | gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10;
   wire 	 pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11) | gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11;
   wire 	 pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12) | gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12;
   wire 	 pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13) | gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13;
   wire 	 pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14) | gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14;
   wire 	 pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15) | gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15;
   wire 	 pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
   wire 	 gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16) | gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16;
   assign Y[0] = pp_0;
   assign Y[1] = pp_1 ^ gg_0;
   assign Y[2] = pp_2 ^ gg_1_gg_0;
   assign Y[3] = pp_3 ^ gg_2_gg_1_gg_0;
   assign Y[4] = pp_4 ^ gg_3_gg_2_gg_1_gg_0;
   assign Y[5] = pp_5 ^ gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[6] = pp_6 ^ gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[7] = pp_7 ^ gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[8] = pp_8 ^ gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[9] = pp_9 ^ gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[10] = pp_10 ^ gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[11] = pp_11 ^ gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[12] = pp_12 ^ gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[13] = pp_13 ^ gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[14] = pp_14 ^ gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[15] = pp_15 ^ gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[16] = pp_16 ^ gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[17] = pp_17 ^ gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[18] = pp_18 ^ gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[19] = pp_19 ^ gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[20] = pp_20 ^ gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[21] = pp_21 ^ gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[22] = pp_22 ^ gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[23] = pp_23 ^ gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[24] = pp_24 ^ gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[25] = pp_25 ^ gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[26] = pp_26 ^ gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[27] = pp_27 ^ gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[28] = pp_28 ^ gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[29] = pp_29 ^ gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[30] = pp_30 ^ gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
   assign Y[31] = pp_31 ^ gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
`endif
endmodule // ppa32


