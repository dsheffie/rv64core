`ifndef __fp_cmp_hdr__
`define __fp_cmp_hdr__

typedef enum logic [3:0] 
{
 CMP_NONE,
 CMP_LT,
 CMP_LE,
 CMP_EQ
} fp_cmp_t;

`endif
