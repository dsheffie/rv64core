`include "machine.vh"

module ppa64(A, B, Y);
input [63:0] A;
input [63:0] B;
output [63:0] Y;
`ifdef FPGA
   assign Y = A+B;
`else   
wire pp_0 = A[0] ^ B[0];
wire gg_0 = A[0] & B[0];
wire pp_1 = A[1] ^ B[1];
wire gg_1 = A[1] & B[1];
wire pp_2 = A[2] ^ B[2];
wire gg_2 = A[2] & B[2];
wire pp_3 = A[3] ^ B[3];
wire gg_3 = A[3] & B[3];
wire pp_4 = A[4] ^ B[4];
wire gg_4 = A[4] & B[4];
wire pp_5 = A[5] ^ B[5];
wire gg_5 = A[5] & B[5];
wire pp_6 = A[6] ^ B[6];
wire gg_6 = A[6] & B[6];
wire pp_7 = A[7] ^ B[7];
wire gg_7 = A[7] & B[7];
wire pp_8 = A[8] ^ B[8];
wire gg_8 = A[8] & B[8];
wire pp_9 = A[9] ^ B[9];
wire gg_9 = A[9] & B[9];
wire pp_10 = A[10] ^ B[10];
wire gg_10 = A[10] & B[10];
wire pp_11 = A[11] ^ B[11];
wire gg_11 = A[11] & B[11];
wire pp_12 = A[12] ^ B[12];
wire gg_12 = A[12] & B[12];
wire pp_13 = A[13] ^ B[13];
wire gg_13 = A[13] & B[13];
wire pp_14 = A[14] ^ B[14];
wire gg_14 = A[14] & B[14];
wire pp_15 = A[15] ^ B[15];
wire gg_15 = A[15] & B[15];
wire pp_16 = A[16] ^ B[16];
wire gg_16 = A[16] & B[16];
wire pp_17 = A[17] ^ B[17];
wire gg_17 = A[17] & B[17];
wire pp_18 = A[18] ^ B[18];
wire gg_18 = A[18] & B[18];
wire pp_19 = A[19] ^ B[19];
wire gg_19 = A[19] & B[19];
wire pp_20 = A[20] ^ B[20];
wire gg_20 = A[20] & B[20];
wire pp_21 = A[21] ^ B[21];
wire gg_21 = A[21] & B[21];
wire pp_22 = A[22] ^ B[22];
wire gg_22 = A[22] & B[22];
wire pp_23 = A[23] ^ B[23];
wire gg_23 = A[23] & B[23];
wire pp_24 = A[24] ^ B[24];
wire gg_24 = A[24] & B[24];
wire pp_25 = A[25] ^ B[25];
wire gg_25 = A[25] & B[25];
wire pp_26 = A[26] ^ B[26];
wire gg_26 = A[26] & B[26];
wire pp_27 = A[27] ^ B[27];
wire gg_27 = A[27] & B[27];
wire pp_28 = A[28] ^ B[28];
wire gg_28 = A[28] & B[28];
wire pp_29 = A[29] ^ B[29];
wire gg_29 = A[29] & B[29];
wire pp_30 = A[30] ^ B[30];
wire gg_30 = A[30] & B[30];
wire pp_31 = A[31] ^ B[31];
wire gg_31 = A[31] & B[31];
wire pp_32 = A[32] ^ B[32];
wire gg_32 = A[32] & B[32];
wire pp_33 = A[33] ^ B[33];
wire gg_33 = A[33] & B[33];
wire pp_34 = A[34] ^ B[34];
wire gg_34 = A[34] & B[34];
wire pp_35 = A[35] ^ B[35];
wire gg_35 = A[35] & B[35];
wire pp_36 = A[36] ^ B[36];
wire gg_36 = A[36] & B[36];
wire pp_37 = A[37] ^ B[37];
wire gg_37 = A[37] & B[37];
wire pp_38 = A[38] ^ B[38];
wire gg_38 = A[38] & B[38];
wire pp_39 = A[39] ^ B[39];
wire gg_39 = A[39] & B[39];
wire pp_40 = A[40] ^ B[40];
wire gg_40 = A[40] & B[40];
wire pp_41 = A[41] ^ B[41];
wire gg_41 = A[41] & B[41];
wire pp_42 = A[42] ^ B[42];
wire gg_42 = A[42] & B[42];
wire pp_43 = A[43] ^ B[43];
wire gg_43 = A[43] & B[43];
wire pp_44 = A[44] ^ B[44];
wire gg_44 = A[44] & B[44];
wire pp_45 = A[45] ^ B[45];
wire gg_45 = A[45] & B[45];
wire pp_46 = A[46] ^ B[46];
wire gg_46 = A[46] & B[46];
wire pp_47 = A[47] ^ B[47];
wire gg_47 = A[47] & B[47];
wire pp_48 = A[48] ^ B[48];
wire gg_48 = A[48] & B[48];
wire pp_49 = A[49] ^ B[49];
wire gg_49 = A[49] & B[49];
wire pp_50 = A[50] ^ B[50];
wire gg_50 = A[50] & B[50];
wire pp_51 = A[51] ^ B[51];
wire gg_51 = A[51] & B[51];
wire pp_52 = A[52] ^ B[52];
wire gg_52 = A[52] & B[52];
wire pp_53 = A[53] ^ B[53];
wire gg_53 = A[53] & B[53];
wire pp_54 = A[54] ^ B[54];
wire gg_54 = A[54] & B[54];
wire pp_55 = A[55] ^ B[55];
wire gg_55 = A[55] & B[55];
wire pp_56 = A[56] ^ B[56];
wire gg_56 = A[56] & B[56];
wire pp_57 = A[57] ^ B[57];
wire gg_57 = A[57] & B[57];
wire pp_58 = A[58] ^ B[58];
wire gg_58 = A[58] & B[58];
wire pp_59 = A[59] ^ B[59];
wire gg_59 = A[59] & B[59];
wire pp_60 = A[60] ^ B[60];
wire gg_60 = A[60] & B[60];
wire pp_61 = A[61] ^ B[61];
wire gg_61 = A[61] & B[61];
wire pp_62 = A[62] ^ B[62];
wire gg_62 = A[62] & B[62];
wire pp_63 = A[63] ^ B[63];
wire gg_63 = A[63] & B[63];
wire pp_1_pp_0 = pp_1 & pp_0;
wire gg_1_gg_0 = (gg_0 & pp_1) | gg_1;
wire pp_2_pp_1 = pp_2 & pp_1;
wire gg_2_gg_1 = (gg_1 & pp_2) | gg_2;
wire pp_3_pp_2 = pp_3 & pp_2;
wire gg_3_gg_2 = (gg_2 & pp_3) | gg_3;
wire pp_4_pp_3 = pp_4 & pp_3;
wire gg_4_gg_3 = (gg_3 & pp_4) | gg_4;
wire pp_5_pp_4 = pp_5 & pp_4;
wire gg_5_gg_4 = (gg_4 & pp_5) | gg_5;
wire pp_6_pp_5 = pp_6 & pp_5;
wire gg_6_gg_5 = (gg_5 & pp_6) | gg_6;
wire pp_7_pp_6 = pp_7 & pp_6;
wire gg_7_gg_6 = (gg_6 & pp_7) | gg_7;
wire pp_8_pp_7 = pp_8 & pp_7;
wire gg_8_gg_7 = (gg_7 & pp_8) | gg_8;
wire pp_9_pp_8 = pp_9 & pp_8;
wire gg_9_gg_8 = (gg_8 & pp_9) | gg_9;
wire pp_10_pp_9 = pp_10 & pp_9;
wire gg_10_gg_9 = (gg_9 & pp_10) | gg_10;
wire pp_11_pp_10 = pp_11 & pp_10;
wire gg_11_gg_10 = (gg_10 & pp_11) | gg_11;
wire pp_12_pp_11 = pp_12 & pp_11;
wire gg_12_gg_11 = (gg_11 & pp_12) | gg_12;
wire pp_13_pp_12 = pp_13 & pp_12;
wire gg_13_gg_12 = (gg_12 & pp_13) | gg_13;
wire pp_14_pp_13 = pp_14 & pp_13;
wire gg_14_gg_13 = (gg_13 & pp_14) | gg_14;
wire pp_15_pp_14 = pp_15 & pp_14;
wire gg_15_gg_14 = (gg_14 & pp_15) | gg_15;
wire pp_16_pp_15 = pp_16 & pp_15;
wire gg_16_gg_15 = (gg_15 & pp_16) | gg_16;
wire pp_17_pp_16 = pp_17 & pp_16;
wire gg_17_gg_16 = (gg_16 & pp_17) | gg_17;
wire pp_18_pp_17 = pp_18 & pp_17;
wire gg_18_gg_17 = (gg_17 & pp_18) | gg_18;
wire pp_19_pp_18 = pp_19 & pp_18;
wire gg_19_gg_18 = (gg_18 & pp_19) | gg_19;
wire pp_20_pp_19 = pp_20 & pp_19;
wire gg_20_gg_19 = (gg_19 & pp_20) | gg_20;
wire pp_21_pp_20 = pp_21 & pp_20;
wire gg_21_gg_20 = (gg_20 & pp_21) | gg_21;
wire pp_22_pp_21 = pp_22 & pp_21;
wire gg_22_gg_21 = (gg_21 & pp_22) | gg_22;
wire pp_23_pp_22 = pp_23 & pp_22;
wire gg_23_gg_22 = (gg_22 & pp_23) | gg_23;
wire pp_24_pp_23 = pp_24 & pp_23;
wire gg_24_gg_23 = (gg_23 & pp_24) | gg_24;
wire pp_25_pp_24 = pp_25 & pp_24;
wire gg_25_gg_24 = (gg_24 & pp_25) | gg_25;
wire pp_26_pp_25 = pp_26 & pp_25;
wire gg_26_gg_25 = (gg_25 & pp_26) | gg_26;
wire pp_27_pp_26 = pp_27 & pp_26;
wire gg_27_gg_26 = (gg_26 & pp_27) | gg_27;
wire pp_28_pp_27 = pp_28 & pp_27;
wire gg_28_gg_27 = (gg_27 & pp_28) | gg_28;
wire pp_29_pp_28 = pp_29 & pp_28;
wire gg_29_gg_28 = (gg_28 & pp_29) | gg_29;
wire pp_30_pp_29 = pp_30 & pp_29;
wire gg_30_gg_29 = (gg_29 & pp_30) | gg_30;
wire pp_31_pp_30 = pp_31 & pp_30;
wire gg_31_gg_30 = (gg_30 & pp_31) | gg_31;
wire pp_32_pp_31 = pp_32 & pp_31;
wire gg_32_gg_31 = (gg_31 & pp_32) | gg_32;
wire pp_33_pp_32 = pp_33 & pp_32;
wire gg_33_gg_32 = (gg_32 & pp_33) | gg_33;
wire pp_34_pp_33 = pp_34 & pp_33;
wire gg_34_gg_33 = (gg_33 & pp_34) | gg_34;
wire pp_35_pp_34 = pp_35 & pp_34;
wire gg_35_gg_34 = (gg_34 & pp_35) | gg_35;
wire pp_36_pp_35 = pp_36 & pp_35;
wire gg_36_gg_35 = (gg_35 & pp_36) | gg_36;
wire pp_37_pp_36 = pp_37 & pp_36;
wire gg_37_gg_36 = (gg_36 & pp_37) | gg_37;
wire pp_38_pp_37 = pp_38 & pp_37;
wire gg_38_gg_37 = (gg_37 & pp_38) | gg_38;
wire pp_39_pp_38 = pp_39 & pp_38;
wire gg_39_gg_38 = (gg_38 & pp_39) | gg_39;
wire pp_40_pp_39 = pp_40 & pp_39;
wire gg_40_gg_39 = (gg_39 & pp_40) | gg_40;
wire pp_41_pp_40 = pp_41 & pp_40;
wire gg_41_gg_40 = (gg_40 & pp_41) | gg_41;
wire pp_42_pp_41 = pp_42 & pp_41;
wire gg_42_gg_41 = (gg_41 & pp_42) | gg_42;
wire pp_43_pp_42 = pp_43 & pp_42;
wire gg_43_gg_42 = (gg_42 & pp_43) | gg_43;
wire pp_44_pp_43 = pp_44 & pp_43;
wire gg_44_gg_43 = (gg_43 & pp_44) | gg_44;
wire pp_45_pp_44 = pp_45 & pp_44;
wire gg_45_gg_44 = (gg_44 & pp_45) | gg_45;
wire pp_46_pp_45 = pp_46 & pp_45;
wire gg_46_gg_45 = (gg_45 & pp_46) | gg_46;
wire pp_47_pp_46 = pp_47 & pp_46;
wire gg_47_gg_46 = (gg_46 & pp_47) | gg_47;
wire pp_48_pp_47 = pp_48 & pp_47;
wire gg_48_gg_47 = (gg_47 & pp_48) | gg_48;
wire pp_49_pp_48 = pp_49 & pp_48;
wire gg_49_gg_48 = (gg_48 & pp_49) | gg_49;
wire pp_50_pp_49 = pp_50 & pp_49;
wire gg_50_gg_49 = (gg_49 & pp_50) | gg_50;
wire pp_51_pp_50 = pp_51 & pp_50;
wire gg_51_gg_50 = (gg_50 & pp_51) | gg_51;
wire pp_52_pp_51 = pp_52 & pp_51;
wire gg_52_gg_51 = (gg_51 & pp_52) | gg_52;
wire pp_53_pp_52 = pp_53 & pp_52;
wire gg_53_gg_52 = (gg_52 & pp_53) | gg_53;
wire pp_54_pp_53 = pp_54 & pp_53;
wire gg_54_gg_53 = (gg_53 & pp_54) | gg_54;
wire pp_55_pp_54 = pp_55 & pp_54;
wire gg_55_gg_54 = (gg_54 & pp_55) | gg_55;
wire pp_56_pp_55 = pp_56 & pp_55;
wire gg_56_gg_55 = (gg_55 & pp_56) | gg_56;
wire pp_57_pp_56 = pp_57 & pp_56;
wire gg_57_gg_56 = (gg_56 & pp_57) | gg_57;
wire pp_58_pp_57 = pp_58 & pp_57;
wire gg_58_gg_57 = (gg_57 & pp_58) | gg_58;
wire pp_59_pp_58 = pp_59 & pp_58;
wire gg_59_gg_58 = (gg_58 & pp_59) | gg_59;
wire pp_60_pp_59 = pp_60 & pp_59;
wire gg_60_gg_59 = (gg_59 & pp_60) | gg_60;
wire pp_61_pp_60 = pp_61 & pp_60;
wire gg_61_gg_60 = (gg_60 & pp_61) | gg_61;
wire pp_62_pp_61 = pp_62 & pp_61;
wire gg_62_gg_61 = (gg_61 & pp_62) | gg_62;
wire pp_63_pp_62 = pp_63 & pp_62;
wire gg_63_gg_62 = (gg_62 & pp_63) | gg_63;
wire pp_2_pp_1_pp_0 = pp_2_pp_1 & pp_0;
wire gg_2_gg_1_gg_0 = (gg_0 & pp_2_pp_1) | gg_2_gg_1;
wire pp_3_pp_2_pp_1_pp_0 = pp_3_pp_2 & pp_1_pp_0;
wire gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_3_pp_2) | gg_3_gg_2;
wire pp_4_pp_3_pp_2_pp_1 = pp_4_pp_3 & pp_2_pp_1;
wire gg_4_gg_3_gg_2_gg_1 = (gg_2_gg_1 & pp_4_pp_3) | gg_4_gg_3;
wire pp_5_pp_4_pp_3_pp_2 = pp_5_pp_4 & pp_3_pp_2;
wire gg_5_gg_4_gg_3_gg_2 = (gg_3_gg_2 & pp_5_pp_4) | gg_5_gg_4;
wire pp_6_pp_5_pp_4_pp_3 = pp_6_pp_5 & pp_4_pp_3;
wire gg_6_gg_5_gg_4_gg_3 = (gg_4_gg_3 & pp_6_pp_5) | gg_6_gg_5;
wire pp_7_pp_6_pp_5_pp_4 = pp_7_pp_6 & pp_5_pp_4;
wire gg_7_gg_6_gg_5_gg_4 = (gg_5_gg_4 & pp_7_pp_6) | gg_7_gg_6;
wire pp_8_pp_7_pp_6_pp_5 = pp_8_pp_7 & pp_6_pp_5;
wire gg_8_gg_7_gg_6_gg_5 = (gg_6_gg_5 & pp_8_pp_7) | gg_8_gg_7;
wire pp_9_pp_8_pp_7_pp_6 = pp_9_pp_8 & pp_7_pp_6;
wire gg_9_gg_8_gg_7_gg_6 = (gg_7_gg_6 & pp_9_pp_8) | gg_9_gg_8;
wire pp_10_pp_9_pp_8_pp_7 = pp_10_pp_9 & pp_8_pp_7;
wire gg_10_gg_9_gg_8_gg_7 = (gg_8_gg_7 & pp_10_pp_9) | gg_10_gg_9;
wire pp_11_pp_10_pp_9_pp_8 = pp_11_pp_10 & pp_9_pp_8;
wire gg_11_gg_10_gg_9_gg_8 = (gg_9_gg_8 & pp_11_pp_10) | gg_11_gg_10;
wire pp_12_pp_11_pp_10_pp_9 = pp_12_pp_11 & pp_10_pp_9;
wire gg_12_gg_11_gg_10_gg_9 = (gg_10_gg_9 & pp_12_pp_11) | gg_12_gg_11;
wire pp_13_pp_12_pp_11_pp_10 = pp_13_pp_12 & pp_11_pp_10;
wire gg_13_gg_12_gg_11_gg_10 = (gg_11_gg_10 & pp_13_pp_12) | gg_13_gg_12;
wire pp_14_pp_13_pp_12_pp_11 = pp_14_pp_13 & pp_12_pp_11;
wire gg_14_gg_13_gg_12_gg_11 = (gg_12_gg_11 & pp_14_pp_13) | gg_14_gg_13;
wire pp_15_pp_14_pp_13_pp_12 = pp_15_pp_14 & pp_13_pp_12;
wire gg_15_gg_14_gg_13_gg_12 = (gg_13_gg_12 & pp_15_pp_14) | gg_15_gg_14;
wire pp_16_pp_15_pp_14_pp_13 = pp_16_pp_15 & pp_14_pp_13;
wire gg_16_gg_15_gg_14_gg_13 = (gg_14_gg_13 & pp_16_pp_15) | gg_16_gg_15;
wire pp_17_pp_16_pp_15_pp_14 = pp_17_pp_16 & pp_15_pp_14;
wire gg_17_gg_16_gg_15_gg_14 = (gg_15_gg_14 & pp_17_pp_16) | gg_17_gg_16;
wire pp_18_pp_17_pp_16_pp_15 = pp_18_pp_17 & pp_16_pp_15;
wire gg_18_gg_17_gg_16_gg_15 = (gg_16_gg_15 & pp_18_pp_17) | gg_18_gg_17;
wire pp_19_pp_18_pp_17_pp_16 = pp_19_pp_18 & pp_17_pp_16;
wire gg_19_gg_18_gg_17_gg_16 = (gg_17_gg_16 & pp_19_pp_18) | gg_19_gg_18;
wire pp_20_pp_19_pp_18_pp_17 = pp_20_pp_19 & pp_18_pp_17;
wire gg_20_gg_19_gg_18_gg_17 = (gg_18_gg_17 & pp_20_pp_19) | gg_20_gg_19;
wire pp_21_pp_20_pp_19_pp_18 = pp_21_pp_20 & pp_19_pp_18;
wire gg_21_gg_20_gg_19_gg_18 = (gg_19_gg_18 & pp_21_pp_20) | gg_21_gg_20;
wire pp_22_pp_21_pp_20_pp_19 = pp_22_pp_21 & pp_20_pp_19;
wire gg_22_gg_21_gg_20_gg_19 = (gg_20_gg_19 & pp_22_pp_21) | gg_22_gg_21;
wire pp_23_pp_22_pp_21_pp_20 = pp_23_pp_22 & pp_21_pp_20;
wire gg_23_gg_22_gg_21_gg_20 = (gg_21_gg_20 & pp_23_pp_22) | gg_23_gg_22;
wire pp_24_pp_23_pp_22_pp_21 = pp_24_pp_23 & pp_22_pp_21;
wire gg_24_gg_23_gg_22_gg_21 = (gg_22_gg_21 & pp_24_pp_23) | gg_24_gg_23;
wire pp_25_pp_24_pp_23_pp_22 = pp_25_pp_24 & pp_23_pp_22;
wire gg_25_gg_24_gg_23_gg_22 = (gg_23_gg_22 & pp_25_pp_24) | gg_25_gg_24;
wire pp_26_pp_25_pp_24_pp_23 = pp_26_pp_25 & pp_24_pp_23;
wire gg_26_gg_25_gg_24_gg_23 = (gg_24_gg_23 & pp_26_pp_25) | gg_26_gg_25;
wire pp_27_pp_26_pp_25_pp_24 = pp_27_pp_26 & pp_25_pp_24;
wire gg_27_gg_26_gg_25_gg_24 = (gg_25_gg_24 & pp_27_pp_26) | gg_27_gg_26;
wire pp_28_pp_27_pp_26_pp_25 = pp_28_pp_27 & pp_26_pp_25;
wire gg_28_gg_27_gg_26_gg_25 = (gg_26_gg_25 & pp_28_pp_27) | gg_28_gg_27;
wire pp_29_pp_28_pp_27_pp_26 = pp_29_pp_28 & pp_27_pp_26;
wire gg_29_gg_28_gg_27_gg_26 = (gg_27_gg_26 & pp_29_pp_28) | gg_29_gg_28;
wire pp_30_pp_29_pp_28_pp_27 = pp_30_pp_29 & pp_28_pp_27;
wire gg_30_gg_29_gg_28_gg_27 = (gg_28_gg_27 & pp_30_pp_29) | gg_30_gg_29;
wire pp_31_pp_30_pp_29_pp_28 = pp_31_pp_30 & pp_29_pp_28;
wire gg_31_gg_30_gg_29_gg_28 = (gg_29_gg_28 & pp_31_pp_30) | gg_31_gg_30;
wire pp_32_pp_31_pp_30_pp_29 = pp_32_pp_31 & pp_30_pp_29;
wire gg_32_gg_31_gg_30_gg_29 = (gg_30_gg_29 & pp_32_pp_31) | gg_32_gg_31;
wire pp_33_pp_32_pp_31_pp_30 = pp_33_pp_32 & pp_31_pp_30;
wire gg_33_gg_32_gg_31_gg_30 = (gg_31_gg_30 & pp_33_pp_32) | gg_33_gg_32;
wire pp_34_pp_33_pp_32_pp_31 = pp_34_pp_33 & pp_32_pp_31;
wire gg_34_gg_33_gg_32_gg_31 = (gg_32_gg_31 & pp_34_pp_33) | gg_34_gg_33;
wire pp_35_pp_34_pp_33_pp_32 = pp_35_pp_34 & pp_33_pp_32;
wire gg_35_gg_34_gg_33_gg_32 = (gg_33_gg_32 & pp_35_pp_34) | gg_35_gg_34;
wire pp_36_pp_35_pp_34_pp_33 = pp_36_pp_35 & pp_34_pp_33;
wire gg_36_gg_35_gg_34_gg_33 = (gg_34_gg_33 & pp_36_pp_35) | gg_36_gg_35;
wire pp_37_pp_36_pp_35_pp_34 = pp_37_pp_36 & pp_35_pp_34;
wire gg_37_gg_36_gg_35_gg_34 = (gg_35_gg_34 & pp_37_pp_36) | gg_37_gg_36;
wire pp_38_pp_37_pp_36_pp_35 = pp_38_pp_37 & pp_36_pp_35;
wire gg_38_gg_37_gg_36_gg_35 = (gg_36_gg_35 & pp_38_pp_37) | gg_38_gg_37;
wire pp_39_pp_38_pp_37_pp_36 = pp_39_pp_38 & pp_37_pp_36;
wire gg_39_gg_38_gg_37_gg_36 = (gg_37_gg_36 & pp_39_pp_38) | gg_39_gg_38;
wire pp_40_pp_39_pp_38_pp_37 = pp_40_pp_39 & pp_38_pp_37;
wire gg_40_gg_39_gg_38_gg_37 = (gg_38_gg_37 & pp_40_pp_39) | gg_40_gg_39;
wire pp_41_pp_40_pp_39_pp_38 = pp_41_pp_40 & pp_39_pp_38;
wire gg_41_gg_40_gg_39_gg_38 = (gg_39_gg_38 & pp_41_pp_40) | gg_41_gg_40;
wire pp_42_pp_41_pp_40_pp_39 = pp_42_pp_41 & pp_40_pp_39;
wire gg_42_gg_41_gg_40_gg_39 = (gg_40_gg_39 & pp_42_pp_41) | gg_42_gg_41;
wire pp_43_pp_42_pp_41_pp_40 = pp_43_pp_42 & pp_41_pp_40;
wire gg_43_gg_42_gg_41_gg_40 = (gg_41_gg_40 & pp_43_pp_42) | gg_43_gg_42;
wire pp_44_pp_43_pp_42_pp_41 = pp_44_pp_43 & pp_42_pp_41;
wire gg_44_gg_43_gg_42_gg_41 = (gg_42_gg_41 & pp_44_pp_43) | gg_44_gg_43;
wire pp_45_pp_44_pp_43_pp_42 = pp_45_pp_44 & pp_43_pp_42;
wire gg_45_gg_44_gg_43_gg_42 = (gg_43_gg_42 & pp_45_pp_44) | gg_45_gg_44;
wire pp_46_pp_45_pp_44_pp_43 = pp_46_pp_45 & pp_44_pp_43;
wire gg_46_gg_45_gg_44_gg_43 = (gg_44_gg_43 & pp_46_pp_45) | gg_46_gg_45;
wire pp_47_pp_46_pp_45_pp_44 = pp_47_pp_46 & pp_45_pp_44;
wire gg_47_gg_46_gg_45_gg_44 = (gg_45_gg_44 & pp_47_pp_46) | gg_47_gg_46;
wire pp_48_pp_47_pp_46_pp_45 = pp_48_pp_47 & pp_46_pp_45;
wire gg_48_gg_47_gg_46_gg_45 = (gg_46_gg_45 & pp_48_pp_47) | gg_48_gg_47;
wire pp_49_pp_48_pp_47_pp_46 = pp_49_pp_48 & pp_47_pp_46;
wire gg_49_gg_48_gg_47_gg_46 = (gg_47_gg_46 & pp_49_pp_48) | gg_49_gg_48;
wire pp_50_pp_49_pp_48_pp_47 = pp_50_pp_49 & pp_48_pp_47;
wire gg_50_gg_49_gg_48_gg_47 = (gg_48_gg_47 & pp_50_pp_49) | gg_50_gg_49;
wire pp_51_pp_50_pp_49_pp_48 = pp_51_pp_50 & pp_49_pp_48;
wire gg_51_gg_50_gg_49_gg_48 = (gg_49_gg_48 & pp_51_pp_50) | gg_51_gg_50;
wire pp_52_pp_51_pp_50_pp_49 = pp_52_pp_51 & pp_50_pp_49;
wire gg_52_gg_51_gg_50_gg_49 = (gg_50_gg_49 & pp_52_pp_51) | gg_52_gg_51;
wire pp_53_pp_52_pp_51_pp_50 = pp_53_pp_52 & pp_51_pp_50;
wire gg_53_gg_52_gg_51_gg_50 = (gg_51_gg_50 & pp_53_pp_52) | gg_53_gg_52;
wire pp_54_pp_53_pp_52_pp_51 = pp_54_pp_53 & pp_52_pp_51;
wire gg_54_gg_53_gg_52_gg_51 = (gg_52_gg_51 & pp_54_pp_53) | gg_54_gg_53;
wire pp_55_pp_54_pp_53_pp_52 = pp_55_pp_54 & pp_53_pp_52;
wire gg_55_gg_54_gg_53_gg_52 = (gg_53_gg_52 & pp_55_pp_54) | gg_55_gg_54;
wire pp_56_pp_55_pp_54_pp_53 = pp_56_pp_55 & pp_54_pp_53;
wire gg_56_gg_55_gg_54_gg_53 = (gg_54_gg_53 & pp_56_pp_55) | gg_56_gg_55;
wire pp_57_pp_56_pp_55_pp_54 = pp_57_pp_56 & pp_55_pp_54;
wire gg_57_gg_56_gg_55_gg_54 = (gg_55_gg_54 & pp_57_pp_56) | gg_57_gg_56;
wire pp_58_pp_57_pp_56_pp_55 = pp_58_pp_57 & pp_56_pp_55;
wire gg_58_gg_57_gg_56_gg_55 = (gg_56_gg_55 & pp_58_pp_57) | gg_58_gg_57;
wire pp_59_pp_58_pp_57_pp_56 = pp_59_pp_58 & pp_57_pp_56;
wire gg_59_gg_58_gg_57_gg_56 = (gg_57_gg_56 & pp_59_pp_58) | gg_59_gg_58;
wire pp_60_pp_59_pp_58_pp_57 = pp_60_pp_59 & pp_58_pp_57;
wire gg_60_gg_59_gg_58_gg_57 = (gg_58_gg_57 & pp_60_pp_59) | gg_60_gg_59;
wire pp_61_pp_60_pp_59_pp_58 = pp_61_pp_60 & pp_59_pp_58;
wire gg_61_gg_60_gg_59_gg_58 = (gg_59_gg_58 & pp_61_pp_60) | gg_61_gg_60;
wire pp_62_pp_61_pp_60_pp_59 = pp_62_pp_61 & pp_60_pp_59;
wire gg_62_gg_61_gg_60_gg_59 = (gg_60_gg_59 & pp_62_pp_61) | gg_62_gg_61;
wire pp_63_pp_62_pp_61_pp_60 = pp_63_pp_62 & pp_61_pp_60;
wire gg_63_gg_62_gg_61_gg_60 = (gg_61_gg_60 & pp_63_pp_62) | gg_63_gg_62;
wire pp_4_pp_3_pp_2_pp_1_pp_0 = pp_4_pp_3_pp_2_pp_1 & pp_0;
wire gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_4_pp_3_pp_2_pp_1) | gg_4_gg_3_gg_2_gg_1;
wire pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
wire gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_5_pp_4_pp_3_pp_2) | gg_5_gg_4_gg_3_gg_2;
wire pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
wire gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_6_pp_5_pp_4_pp_3) | gg_6_gg_5_gg_4_gg_3;
wire pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
wire gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_7_pp_6_pp_5_pp_4) | gg_7_gg_6_gg_5_gg_4;
wire pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 = pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1;
wire gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 = (gg_4_gg_3_gg_2_gg_1 & pp_8_pp_7_pp_6_pp_5) | gg_8_gg_7_gg_6_gg_5;
wire pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 = pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2;
wire gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 = (gg_5_gg_4_gg_3_gg_2 & pp_9_pp_8_pp_7_pp_6) | gg_9_gg_8_gg_7_gg_6;
wire pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 = pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3;
wire gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 = (gg_6_gg_5_gg_4_gg_3 & pp_10_pp_9_pp_8_pp_7) | gg_10_gg_9_gg_8_gg_7;
wire pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 = pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4;
wire gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 = (gg_7_gg_6_gg_5_gg_4 & pp_11_pp_10_pp_9_pp_8) | gg_11_gg_10_gg_9_gg_8;
wire pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 = pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5;
wire gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 = (gg_8_gg_7_gg_6_gg_5 & pp_12_pp_11_pp_10_pp_9) | gg_12_gg_11_gg_10_gg_9;
wire pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 = pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6;
wire gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 = (gg_9_gg_8_gg_7_gg_6 & pp_13_pp_12_pp_11_pp_10) | gg_13_gg_12_gg_11_gg_10;
wire pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 = pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7;
wire gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 = (gg_10_gg_9_gg_8_gg_7 & pp_14_pp_13_pp_12_pp_11) | gg_14_gg_13_gg_12_gg_11;
wire pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 = pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8;
wire gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 = (gg_11_gg_10_gg_9_gg_8 & pp_15_pp_14_pp_13_pp_12) | gg_15_gg_14_gg_13_gg_12;
wire pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 = pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9;
wire gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 = (gg_12_gg_11_gg_10_gg_9 & pp_16_pp_15_pp_14_pp_13) | gg_16_gg_15_gg_14_gg_13;
wire pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 = pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10;
wire gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 = (gg_13_gg_12_gg_11_gg_10 & pp_17_pp_16_pp_15_pp_14) | gg_17_gg_16_gg_15_gg_14;
wire pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 = pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11;
wire gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 = (gg_14_gg_13_gg_12_gg_11 & pp_18_pp_17_pp_16_pp_15) | gg_18_gg_17_gg_16_gg_15;
wire pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 = pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12;
wire gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 = (gg_15_gg_14_gg_13_gg_12 & pp_19_pp_18_pp_17_pp_16) | gg_19_gg_18_gg_17_gg_16;
wire pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 = pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13;
wire gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 = (gg_16_gg_15_gg_14_gg_13 & pp_20_pp_19_pp_18_pp_17) | gg_20_gg_19_gg_18_gg_17;
wire pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 = pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14;
wire gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 = (gg_17_gg_16_gg_15_gg_14 & pp_21_pp_20_pp_19_pp_18) | gg_21_gg_20_gg_19_gg_18;
wire pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 = pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15;
wire gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 = (gg_18_gg_17_gg_16_gg_15 & pp_22_pp_21_pp_20_pp_19) | gg_22_gg_21_gg_20_gg_19;
wire pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 = pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16;
wire gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 = (gg_19_gg_18_gg_17_gg_16 & pp_23_pp_22_pp_21_pp_20) | gg_23_gg_22_gg_21_gg_20;
wire pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 = pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17;
wire gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 = (gg_20_gg_19_gg_18_gg_17 & pp_24_pp_23_pp_22_pp_21) | gg_24_gg_23_gg_22_gg_21;
wire pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 = pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18;
wire gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 = (gg_21_gg_20_gg_19_gg_18 & pp_25_pp_24_pp_23_pp_22) | gg_25_gg_24_gg_23_gg_22;
wire pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 = pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19;
wire gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 = (gg_22_gg_21_gg_20_gg_19 & pp_26_pp_25_pp_24_pp_23) | gg_26_gg_25_gg_24_gg_23;
wire pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 = pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20;
wire gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 = (gg_23_gg_22_gg_21_gg_20 & pp_27_pp_26_pp_25_pp_24) | gg_27_gg_26_gg_25_gg_24;
wire pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 = pp_28_pp_27_pp_26_pp_25 & pp_24_pp_23_pp_22_pp_21;
wire gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 = (gg_24_gg_23_gg_22_gg_21 & pp_28_pp_27_pp_26_pp_25) | gg_28_gg_27_gg_26_gg_25;
wire pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 = pp_29_pp_28_pp_27_pp_26 & pp_25_pp_24_pp_23_pp_22;
wire gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 = (gg_25_gg_24_gg_23_gg_22 & pp_29_pp_28_pp_27_pp_26) | gg_29_gg_28_gg_27_gg_26;
wire pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 = pp_30_pp_29_pp_28_pp_27 & pp_26_pp_25_pp_24_pp_23;
wire gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 = (gg_26_gg_25_gg_24_gg_23 & pp_30_pp_29_pp_28_pp_27) | gg_30_gg_29_gg_28_gg_27;
wire pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 = pp_31_pp_30_pp_29_pp_28 & pp_27_pp_26_pp_25_pp_24;
wire gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 = (gg_27_gg_26_gg_25_gg_24 & pp_31_pp_30_pp_29_pp_28) | gg_31_gg_30_gg_29_gg_28;
wire pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 = pp_32_pp_31_pp_30_pp_29 & pp_28_pp_27_pp_26_pp_25;
wire gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25 = (gg_28_gg_27_gg_26_gg_25 & pp_32_pp_31_pp_30_pp_29) | gg_32_gg_31_gg_30_gg_29;
wire pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 = pp_33_pp_32_pp_31_pp_30 & pp_29_pp_28_pp_27_pp_26;
wire gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26 = (gg_29_gg_28_gg_27_gg_26 & pp_33_pp_32_pp_31_pp_30) | gg_33_gg_32_gg_31_gg_30;
wire pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 = pp_34_pp_33_pp_32_pp_31 & pp_30_pp_29_pp_28_pp_27;
wire gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27 = (gg_30_gg_29_gg_28_gg_27 & pp_34_pp_33_pp_32_pp_31) | gg_34_gg_33_gg_32_gg_31;
wire pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 = pp_35_pp_34_pp_33_pp_32 & pp_31_pp_30_pp_29_pp_28;
wire gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28 = (gg_31_gg_30_gg_29_gg_28 & pp_35_pp_34_pp_33_pp_32) | gg_35_gg_34_gg_33_gg_32;
wire pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 = pp_36_pp_35_pp_34_pp_33 & pp_32_pp_31_pp_30_pp_29;
wire gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29 = (gg_32_gg_31_gg_30_gg_29 & pp_36_pp_35_pp_34_pp_33) | gg_36_gg_35_gg_34_gg_33;
wire pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 = pp_37_pp_36_pp_35_pp_34 & pp_33_pp_32_pp_31_pp_30;
wire gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30 = (gg_33_gg_32_gg_31_gg_30 & pp_37_pp_36_pp_35_pp_34) | gg_37_gg_36_gg_35_gg_34;
wire pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 = pp_38_pp_37_pp_36_pp_35 & pp_34_pp_33_pp_32_pp_31;
wire gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31 = (gg_34_gg_33_gg_32_gg_31 & pp_38_pp_37_pp_36_pp_35) | gg_38_gg_37_gg_36_gg_35;
wire pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 = pp_39_pp_38_pp_37_pp_36 & pp_35_pp_34_pp_33_pp_32;
wire gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32 = (gg_35_gg_34_gg_33_gg_32 & pp_39_pp_38_pp_37_pp_36) | gg_39_gg_38_gg_37_gg_36;
wire pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33 = pp_40_pp_39_pp_38_pp_37 & pp_36_pp_35_pp_34_pp_33;
wire gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33 = (gg_36_gg_35_gg_34_gg_33 & pp_40_pp_39_pp_38_pp_37) | gg_40_gg_39_gg_38_gg_37;
wire pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34 = pp_41_pp_40_pp_39_pp_38 & pp_37_pp_36_pp_35_pp_34;
wire gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34 = (gg_37_gg_36_gg_35_gg_34 & pp_41_pp_40_pp_39_pp_38) | gg_41_gg_40_gg_39_gg_38;
wire pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35 = pp_42_pp_41_pp_40_pp_39 & pp_38_pp_37_pp_36_pp_35;
wire gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35 = (gg_38_gg_37_gg_36_gg_35 & pp_42_pp_41_pp_40_pp_39) | gg_42_gg_41_gg_40_gg_39;
wire pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36 = pp_43_pp_42_pp_41_pp_40 & pp_39_pp_38_pp_37_pp_36;
wire gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36 = (gg_39_gg_38_gg_37_gg_36 & pp_43_pp_42_pp_41_pp_40) | gg_43_gg_42_gg_41_gg_40;
wire pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37 = pp_44_pp_43_pp_42_pp_41 & pp_40_pp_39_pp_38_pp_37;
wire gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37 = (gg_40_gg_39_gg_38_gg_37 & pp_44_pp_43_pp_42_pp_41) | gg_44_gg_43_gg_42_gg_41;
wire pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38 = pp_45_pp_44_pp_43_pp_42 & pp_41_pp_40_pp_39_pp_38;
wire gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38 = (gg_41_gg_40_gg_39_gg_38 & pp_45_pp_44_pp_43_pp_42) | gg_45_gg_44_gg_43_gg_42;
wire pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39 = pp_46_pp_45_pp_44_pp_43 & pp_42_pp_41_pp_40_pp_39;
wire gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39 = (gg_42_gg_41_gg_40_gg_39 & pp_46_pp_45_pp_44_pp_43) | gg_46_gg_45_gg_44_gg_43;
wire pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40 = pp_47_pp_46_pp_45_pp_44 & pp_43_pp_42_pp_41_pp_40;
wire gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40 = (gg_43_gg_42_gg_41_gg_40 & pp_47_pp_46_pp_45_pp_44) | gg_47_gg_46_gg_45_gg_44;
wire pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41 = pp_48_pp_47_pp_46_pp_45 & pp_44_pp_43_pp_42_pp_41;
wire gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41 = (gg_44_gg_43_gg_42_gg_41 & pp_48_pp_47_pp_46_pp_45) | gg_48_gg_47_gg_46_gg_45;
wire pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42 = pp_49_pp_48_pp_47_pp_46 & pp_45_pp_44_pp_43_pp_42;
wire gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42 = (gg_45_gg_44_gg_43_gg_42 & pp_49_pp_48_pp_47_pp_46) | gg_49_gg_48_gg_47_gg_46;
wire pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43 = pp_50_pp_49_pp_48_pp_47 & pp_46_pp_45_pp_44_pp_43;
wire gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43 = (gg_46_gg_45_gg_44_gg_43 & pp_50_pp_49_pp_48_pp_47) | gg_50_gg_49_gg_48_gg_47;
wire pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44 = pp_51_pp_50_pp_49_pp_48 & pp_47_pp_46_pp_45_pp_44;
wire gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44 = (gg_47_gg_46_gg_45_gg_44 & pp_51_pp_50_pp_49_pp_48) | gg_51_gg_50_gg_49_gg_48;
wire pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45 = pp_52_pp_51_pp_50_pp_49 & pp_48_pp_47_pp_46_pp_45;
wire gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45 = (gg_48_gg_47_gg_46_gg_45 & pp_52_pp_51_pp_50_pp_49) | gg_52_gg_51_gg_50_gg_49;
wire pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46 = pp_53_pp_52_pp_51_pp_50 & pp_49_pp_48_pp_47_pp_46;
wire gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46 = (gg_49_gg_48_gg_47_gg_46 & pp_53_pp_52_pp_51_pp_50) | gg_53_gg_52_gg_51_gg_50;
wire pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47 = pp_54_pp_53_pp_52_pp_51 & pp_50_pp_49_pp_48_pp_47;
wire gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47 = (gg_50_gg_49_gg_48_gg_47 & pp_54_pp_53_pp_52_pp_51) | gg_54_gg_53_gg_52_gg_51;
wire pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48 = pp_55_pp_54_pp_53_pp_52 & pp_51_pp_50_pp_49_pp_48;
wire gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48 = (gg_51_gg_50_gg_49_gg_48 & pp_55_pp_54_pp_53_pp_52) | gg_55_gg_54_gg_53_gg_52;
wire pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49 = pp_56_pp_55_pp_54_pp_53 & pp_52_pp_51_pp_50_pp_49;
wire gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49 = (gg_52_gg_51_gg_50_gg_49 & pp_56_pp_55_pp_54_pp_53) | gg_56_gg_55_gg_54_gg_53;
wire pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50 = pp_57_pp_56_pp_55_pp_54 & pp_53_pp_52_pp_51_pp_50;
wire gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50 = (gg_53_gg_52_gg_51_gg_50 & pp_57_pp_56_pp_55_pp_54) | gg_57_gg_56_gg_55_gg_54;
wire pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51 = pp_58_pp_57_pp_56_pp_55 & pp_54_pp_53_pp_52_pp_51;
wire gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51 = (gg_54_gg_53_gg_52_gg_51 & pp_58_pp_57_pp_56_pp_55) | gg_58_gg_57_gg_56_gg_55;
wire pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52 = pp_59_pp_58_pp_57_pp_56 & pp_55_pp_54_pp_53_pp_52;
wire gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52 = (gg_55_gg_54_gg_53_gg_52 & pp_59_pp_58_pp_57_pp_56) | gg_59_gg_58_gg_57_gg_56;
wire pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53 = pp_60_pp_59_pp_58_pp_57 & pp_56_pp_55_pp_54_pp_53;
wire gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53 = (gg_56_gg_55_gg_54_gg_53 & pp_60_pp_59_pp_58_pp_57) | gg_60_gg_59_gg_58_gg_57;
wire pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54 = pp_61_pp_60_pp_59_pp_58 & pp_57_pp_56_pp_55_pp_54;
wire gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54 = (gg_57_gg_56_gg_55_gg_54 & pp_61_pp_60_pp_59_pp_58) | gg_61_gg_60_gg_59_gg_58;
wire pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55 = pp_62_pp_61_pp_60_pp_59 & pp_58_pp_57_pp_56_pp_55;
wire gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55 = (gg_58_gg_57_gg_56_gg_55 & pp_62_pp_61_pp_60_pp_59) | gg_62_gg_61_gg_60_gg_59;
wire pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56 = pp_63_pp_62_pp_61_pp_60 & pp_59_pp_58_pp_57_pp_56;
wire gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56 = (gg_59_gg_58_gg_57_gg_56 & pp_63_pp_62_pp_61_pp_60) | gg_63_gg_62_gg_61_gg_60;
wire pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 & pp_0;
wire gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1) | gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1;
wire pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
wire gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2) | gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2;
wire pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
wire gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3) | gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3;
wire pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
wire gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4) | gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4;
wire pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_4_gg_3_gg_2_gg_1_gg_0 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5) | gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5;
wire pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6) | gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6;
wire pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7) | gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7;
wire pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8) | gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8;
wire pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 = pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1;
wire gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 = (gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9) | gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9;
wire pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 = pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2;
wire gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 = (gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10) | gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10;
wire pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 = pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3;
wire gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 = (gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11) | gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11;
wire pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 = pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4;
wire gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 = (gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12) | gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12;
wire pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 = pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5;
wire gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 = (gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13) | gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13;
wire pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 = pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6;
wire gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 = (gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14) | gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14;
wire pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 = pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7;
wire gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 = (gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15) | gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15;
wire pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 = pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8;
wire gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 = (gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16) | gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16;
wire pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 = pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9;
wire gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 = (gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17) | gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17;
wire pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 = pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10;
wire gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 = (gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18) | gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18;
wire pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 = pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11;
wire gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 = (gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19) | gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19;
wire pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 = pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12;
wire gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 = (gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20) | gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20;
wire pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 = pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13;
wire gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 = (gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21) | gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21;
wire pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 = pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14;
wire gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 = (gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22) | gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22;
wire pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 = pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15;
wire gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 = (gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23) | gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23;
wire pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 = pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16;
wire gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 = (gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24) | gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24;
wire pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 = pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17;
wire gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 = (gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 & pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25) | gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25;
wire pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 = pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18;
wire gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 = (gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 & pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26) | gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26;
wire pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 = pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19;
wire gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 = (gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 & pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27) | gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27;
wire pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 = pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20;
wire gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 = (gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 & pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28) | gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28;
wire pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 = pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21;
wire gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 = (gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 & pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29) | gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29;
wire pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 = pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22;
wire gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 = (gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 & pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30) | gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30;
wire pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 = pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23;
wire gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 = (gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 & pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31) | gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31;
wire pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 = pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24;
wire gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 = (gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 & pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32) | gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32;
wire pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 = pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33 & pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25;
wire gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25 = (gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25 & pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33) | gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33;
wire pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 = pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34 & pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26;
wire gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26 = (gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26 & pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34) | gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34;
wire pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 = pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35 & pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27;
wire gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27 = (gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27 & pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35) | gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35;
wire pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 = pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36 & pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28;
wire gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28 = (gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28 & pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36) | gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36;
wire pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 = pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37 & pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29;
wire gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29 = (gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29 & pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37) | gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37;
wire pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 = pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38 & pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30;
wire gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30 = (gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30 & pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38) | gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38;
wire pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 = pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39 & pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31;
wire gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31 = (gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31 & pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39) | gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39;
wire pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 = pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40 & pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32;
wire gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32 = (gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32 & pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40) | gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40;
wire pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33 = pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41 & pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33;
wire gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33 = (gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33 & pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41) | gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41;
wire pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34 = pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42 & pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34;
wire gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34 = (gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34 & pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42) | gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42;
wire pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35 = pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43 & pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35;
wire gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35 = (gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35 & pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43) | gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43;
wire pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36 = pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44 & pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36;
wire gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36 = (gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36 & pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44) | gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44;
wire pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37 = pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45 & pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37;
wire gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37 = (gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37 & pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45) | gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45;
wire pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38 = pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46 & pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38;
wire gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38 = (gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38 & pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46) | gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46;
wire pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39 = pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47 & pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39;
wire gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39 = (gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39 & pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47) | gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47;
wire pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40 = pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48 & pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40;
wire gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40 = (gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40 & pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48) | gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48;
wire pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41 = pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49 & pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41;
wire gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41 = (gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41 & pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49) | gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49;
wire pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42 = pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50 & pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42;
wire gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42 = (gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42 & pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50) | gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50;
wire pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43 = pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51 & pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43;
wire gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43 = (gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43 & pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51) | gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51;
wire pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44 = pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52 & pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44;
wire gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44 = (gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44 & pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52) | gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52;
wire pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45 = pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53 & pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45;
wire gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45 = (gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45 & pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53) | gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53;
wire pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46 = pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54 & pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46;
wire gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46 = (gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46 & pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54) | gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54;
wire pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47 = pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55 & pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47;
wire gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47 = (gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47 & pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55) | gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55;
wire pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48 = pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56 & pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48;
wire gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48 = (gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48 & pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56) | gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56;
wire pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 & pp_0;
wire gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1) | gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1;
wire pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
wire gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2) | gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2;
wire pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
wire gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3) | gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3;
wire pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
wire gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4) | gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4;
wire pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_4_gg_3_gg_2_gg_1_gg_0 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5) | gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5;
wire pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6) | gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6;
wire pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7) | gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7;
wire pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8) | gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8;
wire pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9) | gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9;
wire pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10) | gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10;
wire pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11) | gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11;
wire pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12) | gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12;
wire pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13) | gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13;
wire pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14) | gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14;
wire pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15) | gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15;
wire pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16) | gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16;
wire pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 = pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1;
wire gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 = (gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1 & pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17) | gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17;
wire pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 = pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2;
wire gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 = (gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2 & pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18) | gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18;
wire pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 = pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3;
wire gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 = (gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3 & pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19) | gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19;
wire pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 = pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4;
wire gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 = (gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4 & pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20) | gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20;
wire pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 = pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5;
wire gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 = (gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5 & pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21) | gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21;
wire pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 = pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6;
wire gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 = (gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6 & pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22) | gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22;
wire pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 = pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7;
wire gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 = (gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7 & pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23) | gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23;
wire pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 = pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8;
wire gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 = (gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8 & pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24) | gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24;
wire pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 = pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9;
wire gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 = (gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9 & pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25) | gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25;
wire pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 = pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10;
wire gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 = (gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10 & pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26) | gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26;
wire pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 = pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11;
wire gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 = (gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11 & pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27) | gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27;
wire pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 = pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12;
wire gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 = (gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12 & pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28) | gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28;
wire pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 = pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13;
wire gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 = (gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13 & pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29) | gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29;
wire pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 = pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14;
wire gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 = (gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14 & pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30) | gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30;
wire pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 = pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15;
wire gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 = (gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15 & pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31) | gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31;
wire pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 = pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16;
wire gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 = (gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16 & pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32) | gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32;
wire pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 = pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33 & pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17;
wire gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 = (gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17 & pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33) | gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33;
wire pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 = pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34 & pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18;
wire gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 = (gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18 & pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34) | gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34;
wire pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 = pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35 & pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19;
wire gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 = (gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19 & pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35) | gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35;
wire pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 = pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36 & pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20;
wire gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 = (gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20 & pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36) | gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36;
wire pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 = pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37 & pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21;
wire gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 = (gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21 & pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37) | gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37;
wire pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 = pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38 & pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22;
wire gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 = (gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22 & pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38) | gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38;
wire pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 = pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39 & pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23;
wire gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 = (gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23 & pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39) | gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39;
wire pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 = pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40 & pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24;
wire gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 = (gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24 & pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40) | gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40;
wire pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 = pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41 & pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25;
wire gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25 = (gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25 & pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41) | gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41;
wire pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 = pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42 & pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26;
wire gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26 = (gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26 & pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42) | gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42;
wire pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 = pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43 & pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27;
wire gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27 = (gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27 & pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43) | gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43;
wire pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 = pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44 & pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28;
wire gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28 = (gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28 & pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44) | gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44;
wire pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 = pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45 & pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29;
wire gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29 = (gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29 & pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45) | gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45;
wire pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 = pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46 & pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30;
wire gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30 = (gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30 & pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46) | gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46;
wire pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 = pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47 & pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31;
wire gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31 = (gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31 & pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47) | gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47;
wire pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 = pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48 & pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32;
wire gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32 = (gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32 & pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48) | gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48;
wire pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1 & pp_0;
wire gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_0 & pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1) | gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1;
wire pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2 & pp_1_pp_0;
wire gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_1_gg_0 & pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2) | gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2;
wire pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3 & pp_2_pp_1_pp_0;
wire gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_2_gg_1_gg_0 & pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3) | gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3;
wire pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4 & pp_3_pp_2_pp_1_pp_0;
wire gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_3_gg_2_gg_1_gg_0 & pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4) | gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4;
wire pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5 & pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_4_gg_3_gg_2_gg_1_gg_0 & pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5) | gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5;
wire pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6 & pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6) | gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6;
wire pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7 & pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7) | gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7;
wire pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8 & pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8) | gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8;
wire pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9 & pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9) | gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9;
wire pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10 & pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10) | gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10;
wire pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11 & pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11) | gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11;
wire pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12 & pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12) | gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12;
wire pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13 & pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13) | gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13;
wire pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14 & pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14) | gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14;
wire pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15 & pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15) | gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15;
wire pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16 & pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16) | gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16;
wire pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17 & pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17) | gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17;
wire pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18 & pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18) | gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18;
wire pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19 & pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19) | gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19;
wire pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20 & pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20) | gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20;
wire pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21 & pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21) | gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21;
wire pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22 & pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22) | gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22;
wire pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23 & pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23) | gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23;
wire pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24 & pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24) | gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24;
wire pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25 & pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25) | gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25;
wire pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26 & pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26) | gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26;
wire pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27 & pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27) | gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27;
wire pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28 & pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28) | gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28;
wire pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29 & pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29) | gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29;
wire pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30 & pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30) | gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30;
wire pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31 & pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31) | gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31;
wire pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32_pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0 = pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32 & pp_31_pp_30_pp_29_pp_28_pp_27_pp_26_pp_25_pp_24_pp_23_pp_22_pp_21_pp_20_pp_19_pp_18_pp_17_pp_16_pp_15_pp_14_pp_13_pp_12_pp_11_pp_10_pp_9_pp_8_pp_7_pp_6_pp_5_pp_4_pp_3_pp_2_pp_1_pp_0;
wire gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 = (gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0 & pp_63_pp_62_pp_61_pp_60_pp_59_pp_58_pp_57_pp_56_pp_55_pp_54_pp_53_pp_52_pp_51_pp_50_pp_49_pp_48_pp_47_pp_46_pp_45_pp_44_pp_43_pp_42_pp_41_pp_40_pp_39_pp_38_pp_37_pp_36_pp_35_pp_34_pp_33_pp_32) | gg_63_gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32;
assign Y[0] = pp_0;
assign Y[1] = pp_1 ^ gg_0;
assign Y[2] = pp_2 ^ gg_1_gg_0;
assign Y[3] = pp_3 ^ gg_2_gg_1_gg_0;
assign Y[4] = pp_4 ^ gg_3_gg_2_gg_1_gg_0;
assign Y[5] = pp_5 ^ gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[6] = pp_6 ^ gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[7] = pp_7 ^ gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[8] = pp_8 ^ gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[9] = pp_9 ^ gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[10] = pp_10 ^ gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[11] = pp_11 ^ gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[12] = pp_12 ^ gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[13] = pp_13 ^ gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[14] = pp_14 ^ gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[15] = pp_15 ^ gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[16] = pp_16 ^ gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[17] = pp_17 ^ gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[18] = pp_18 ^ gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[19] = pp_19 ^ gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[20] = pp_20 ^ gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[21] = pp_21 ^ gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[22] = pp_22 ^ gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[23] = pp_23 ^ gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[24] = pp_24 ^ gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[25] = pp_25 ^ gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[26] = pp_26 ^ gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[27] = pp_27 ^ gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[28] = pp_28 ^ gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[29] = pp_29 ^ gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[30] = pp_30 ^ gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[31] = pp_31 ^ gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[32] = pp_32 ^ gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[33] = pp_33 ^ gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[34] = pp_34 ^ gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[35] = pp_35 ^ gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[36] = pp_36 ^ gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[37] = pp_37 ^ gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[38] = pp_38 ^ gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[39] = pp_39 ^ gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[40] = pp_40 ^ gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[41] = pp_41 ^ gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[42] = pp_42 ^ gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[43] = pp_43 ^ gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[44] = pp_44 ^ gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[45] = pp_45 ^ gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[46] = pp_46 ^ gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[47] = pp_47 ^ gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[48] = pp_48 ^ gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[49] = pp_49 ^ gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[50] = pp_50 ^ gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[51] = pp_51 ^ gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[52] = pp_52 ^ gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[53] = pp_53 ^ gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[54] = pp_54 ^ gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[55] = pp_55 ^ gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[56] = pp_56 ^ gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[57] = pp_57 ^ gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[58] = pp_58 ^ gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[59] = pp_59 ^ gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[60] = pp_60 ^ gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[61] = pp_61 ^ gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[62] = pp_62 ^ gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
assign Y[63] = pp_63 ^ gg_62_gg_61_gg_60_gg_59_gg_58_gg_57_gg_56_gg_55_gg_54_gg_53_gg_52_gg_51_gg_50_gg_49_gg_48_gg_47_gg_46_gg_45_gg_44_gg_43_gg_42_gg_41_gg_40_gg_39_gg_38_gg_37_gg_36_gg_35_gg_34_gg_33_gg_32_gg_31_gg_30_gg_29_gg_28_gg_27_gg_26_gg_25_gg_24_gg_23_gg_22_gg_21_gg_20_gg_19_gg_18_gg_17_gg_16_gg_15_gg_14_gg_13_gg_12_gg_11_gg_10_gg_9_gg_8_gg_7_gg_6_gg_5_gg_4_gg_3_gg_2_gg_1_gg_0;
`endif // !`ifdef FPGA   
endmodule // ppa64





