module ctz64(A, Y);
input logic [63:0] A;
output logic [6:0] Y;
always_comb
begin
  Y = 'd0;
  casez(A)
   64'b0000000000000000000000000000000000000000000000000000000000000000: Y = 'd64;
   64'b1000000000000000000000000000000000000000000000000000000000000000: Y = 'd63;
   64'b?100000000000000000000000000000000000000000000000000000000000000: Y = 'd62;
   64'b??10000000000000000000000000000000000000000000000000000000000000: Y = 'd61;
   64'b???1000000000000000000000000000000000000000000000000000000000000: Y = 'd60;
   64'b????100000000000000000000000000000000000000000000000000000000000: Y = 'd59;
   64'b?????10000000000000000000000000000000000000000000000000000000000: Y = 'd58;
   64'b??????1000000000000000000000000000000000000000000000000000000000: Y = 'd57;
   64'b???????100000000000000000000000000000000000000000000000000000000: Y = 'd56;
   64'b????????10000000000000000000000000000000000000000000000000000000: Y = 'd55;
   64'b?????????1000000000000000000000000000000000000000000000000000000: Y = 'd54;
   64'b??????????100000000000000000000000000000000000000000000000000000: Y = 'd53;
   64'b???????????10000000000000000000000000000000000000000000000000000: Y = 'd52;
   64'b????????????1000000000000000000000000000000000000000000000000000: Y = 'd51;
   64'b?????????????100000000000000000000000000000000000000000000000000: Y = 'd50;
   64'b??????????????10000000000000000000000000000000000000000000000000: Y = 'd49;
   64'b???????????????1000000000000000000000000000000000000000000000000: Y = 'd48;
   64'b????????????????100000000000000000000000000000000000000000000000: Y = 'd47;
   64'b?????????????????10000000000000000000000000000000000000000000000: Y = 'd46;
   64'b??????????????????1000000000000000000000000000000000000000000000: Y = 'd45;
   64'b???????????????????100000000000000000000000000000000000000000000: Y = 'd44;
   64'b????????????????????10000000000000000000000000000000000000000000: Y = 'd43;
   64'b?????????????????????1000000000000000000000000000000000000000000: Y = 'd42;
   64'b??????????????????????100000000000000000000000000000000000000000: Y = 'd41;
   64'b???????????????????????10000000000000000000000000000000000000000: Y = 'd40;
   64'b????????????????????????1000000000000000000000000000000000000000: Y = 'd39;
   64'b?????????????????????????100000000000000000000000000000000000000: Y = 'd38;
   64'b??????????????????????????10000000000000000000000000000000000000: Y = 'd37;
   64'b???????????????????????????1000000000000000000000000000000000000: Y = 'd36;
   64'b????????????????????????????100000000000000000000000000000000000: Y = 'd35;
   64'b?????????????????????????????10000000000000000000000000000000000: Y = 'd34;
   64'b??????????????????????????????1000000000000000000000000000000000: Y = 'd33;
   64'b???????????????????????????????100000000000000000000000000000000: Y = 'd32;
   64'b????????????????????????????????10000000000000000000000000000000: Y = 'd31;
   64'b?????????????????????????????????1000000000000000000000000000000: Y = 'd30;
   64'b??????????????????????????????????100000000000000000000000000000: Y = 'd29;
   64'b???????????????????????????????????10000000000000000000000000000: Y = 'd28;
   64'b????????????????????????????????????1000000000000000000000000000: Y = 'd27;
   64'b?????????????????????????????????????100000000000000000000000000: Y = 'd26;
   64'b??????????????????????????????????????10000000000000000000000000: Y = 'd25;
   64'b???????????????????????????????????????1000000000000000000000000: Y = 'd24;
   64'b????????????????????????????????????????100000000000000000000000: Y = 'd23;
   64'b?????????????????????????????????????????10000000000000000000000: Y = 'd22;
   64'b??????????????????????????????????????????1000000000000000000000: Y = 'd21;
   64'b???????????????????????????????????????????100000000000000000000: Y = 'd20;
   64'b????????????????????????????????????????????10000000000000000000: Y = 'd19;
   64'b?????????????????????????????????????????????1000000000000000000: Y = 'd18;
   64'b??????????????????????????????????????????????100000000000000000: Y = 'd17;
   64'b???????????????????????????????????????????????10000000000000000: Y = 'd16;
   64'b????????????????????????????????????????????????1000000000000000: Y = 'd15;
   64'b?????????????????????????????????????????????????100000000000000: Y = 'd14;
   64'b??????????????????????????????????????????????????10000000000000: Y = 'd13;
   64'b???????????????????????????????????????????????????1000000000000: Y = 'd12;
   64'b????????????????????????????????????????????????????100000000000: Y = 'd11;
   64'b?????????????????????????????????????????????????????10000000000: Y = 'd10;
   64'b??????????????????????????????????????????????????????1000000000: Y = 'd9;
   64'b???????????????????????????????????????????????????????100000000: Y = 'd8;
   64'b????????????????????????????????????????????????????????10000000: Y = 'd7;
   64'b?????????????????????????????????????????????????????????1000000: Y = 'd6;
   64'b??????????????????????????????????????????????????????????100000: Y = 'd5;
   64'b???????????????????????????????????????????????????????????10000: Y = 'd4;
   64'b????????????????????????????????????????????????????????????1000: Y = 'd3;
   64'b?????????????????????????????????????????????????????????????100: Y = 'd2;
   64'b??????????????????????????????????????????????????????????????10: Y = 'd1;
  default:
    begin
    end
  endcase
end
endmodule
