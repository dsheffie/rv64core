module clz64(A, Y);
input logic [63:0] A;
output logic [6:0] Y;
always_comb
begin
  Y = 'd0;
  casez(A)
    64'b0000000000000000000000000000000000000000000000000000000000000000: Y = 'd64;
    64'b0000000000000000000000000000000000000000000000000000000000000001: Y = 'd63;
    64'b000000000000000000000000000000000000000000000000000000000000001?: Y = 'd62;
    64'b00000000000000000000000000000000000000000000000000000000000001??: Y = 'd61;
    64'b0000000000000000000000000000000000000000000000000000000000001???: Y = 'd60;
    64'b000000000000000000000000000000000000000000000000000000000001????: Y = 'd59;
    64'b00000000000000000000000000000000000000000000000000000000001?????: Y = 'd58;
    64'b0000000000000000000000000000000000000000000000000000000001??????: Y = 'd57;
    64'b000000000000000000000000000000000000000000000000000000001???????: Y = 'd56;
    64'b00000000000000000000000000000000000000000000000000000001????????: Y = 'd55;
    64'b0000000000000000000000000000000000000000000000000000001?????????: Y = 'd54;
    64'b000000000000000000000000000000000000000000000000000001??????????: Y = 'd53;
    64'b00000000000000000000000000000000000000000000000000001???????????: Y = 'd52;
    64'b0000000000000000000000000000000000000000000000000001????????????: Y = 'd51;
    64'b000000000000000000000000000000000000000000000000001?????????????: Y = 'd50;
    64'b00000000000000000000000000000000000000000000000001??????????????: Y = 'd49;
    64'b0000000000000000000000000000000000000000000000001???????????????: Y = 'd48;
    64'b000000000000000000000000000000000000000000000001????????????????: Y = 'd47;
    64'b00000000000000000000000000000000000000000000001?????????????????: Y = 'd46;
    64'b0000000000000000000000000000000000000000000001??????????????????: Y = 'd45;
    64'b000000000000000000000000000000000000000000001???????????????????: Y = 'd44;
    64'b00000000000000000000000000000000000000000001????????????????????: Y = 'd43;
    64'b0000000000000000000000000000000000000000001?????????????????????: Y = 'd42;
    64'b000000000000000000000000000000000000000001??????????????????????: Y = 'd41;
    64'b00000000000000000000000000000000000000001???????????????????????: Y = 'd40;
    64'b0000000000000000000000000000000000000001????????????????????????: Y = 'd39;
    64'b000000000000000000000000000000000000001?????????????????????????: Y = 'd38;
    64'b00000000000000000000000000000000000001??????????????????????????: Y = 'd37;
    64'b0000000000000000000000000000000000001???????????????????????????: Y = 'd36;
    64'b000000000000000000000000000000000001????????????????????????????: Y = 'd35;
    64'b00000000000000000000000000000000001?????????????????????????????: Y = 'd34;
    64'b0000000000000000000000000000000001??????????????????????????????: Y = 'd33;
    64'b000000000000000000000000000000001???????????????????????????????: Y = 'd32;
    64'b00000000000000000000000000000001????????????????????????????????: Y = 'd31;
    64'b0000000000000000000000000000001?????????????????????????????????: Y = 'd30;
    64'b000000000000000000000000000001??????????????????????????????????: Y = 'd29;
    64'b00000000000000000000000000001???????????????????????????????????: Y = 'd28;
    64'b0000000000000000000000000001????????????????????????????????????: Y = 'd27;
    64'b000000000000000000000000001?????????????????????????????????????: Y = 'd26;
    64'b00000000000000000000000001??????????????????????????????????????: Y = 'd25;
    64'b0000000000000000000000001???????????????????????????????????????: Y = 'd24;
    64'b000000000000000000000001????????????????????????????????????????: Y = 'd23;
    64'b00000000000000000000001?????????????????????????????????????????: Y = 'd22;
    64'b0000000000000000000001??????????????????????????????????????????: Y = 'd21;
    64'b000000000000000000001???????????????????????????????????????????: Y = 'd20;
    64'b00000000000000000001????????????????????????????????????????????: Y = 'd19;
    64'b0000000000000000001?????????????????????????????????????????????: Y = 'd18;
    64'b000000000000000001??????????????????????????????????????????????: Y = 'd17;
    64'b00000000000000001???????????????????????????????????????????????: Y = 'd16;
    64'b0000000000000001????????????????????????????????????????????????: Y = 'd15;
    64'b000000000000001?????????????????????????????????????????????????: Y = 'd14;
    64'b00000000000001??????????????????????????????????????????????????: Y = 'd13;
    64'b0000000000001???????????????????????????????????????????????????: Y = 'd12;
    64'b000000000001????????????????????????????????????????????????????: Y = 'd11;
    64'b00000000001?????????????????????????????????????????????????????: Y = 'd10;
    64'b0000000001??????????????????????????????????????????????????????: Y = 'd9;
    64'b000000001???????????????????????????????????????????????????????: Y = 'd8;
    64'b00000001????????????????????????????????????????????????????????: Y = 'd7;
    64'b0000001?????????????????????????????????????????????????????????: Y = 'd6;
    64'b000001??????????????????????????????????????????????????????????: Y = 'd5;
    64'b00001???????????????????????????????????????????????????????????: Y = 'd4;
    64'b0001????????????????????????????????????????????????????????????: Y = 'd3;
    64'b001?????????????????????????????????????????????????????????????: Y = 'd2;
    64'b01??????????????????????????????????????????????????????????????: Y = 'd1;
  default:
    begin
    end
  endcase
end
endmodule
